// Code your design here
`timescale 1ns/1ps


module full_adder(input a,
                  input b,
                  input c,
                  output sum,
                  output carry);
  assign {carry,sum} = a+b+c;
endmodule



module ripple_carry_adder(
  input [3:0]a,
  input [3:0]b,
  input c,
  output [3:0]sum,
  output carry);
  
  wire c1,c2,c3;
  
  full_adder F0(a[0],b[0],c,sum[0],c1);
  full_adder F1(a[1],b[1],c1,sum[1],c2);
  full_adder F2(a[2],b[2],c2,sum[2],c3);
  full_adder F3(a[3],b[3],c3,sum[3],carry);
endmodule
  
