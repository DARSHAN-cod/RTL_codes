// Code your design here
module dff_enable (
    input  wire clk,
    input  wire rst,   
    input  wire en,      
    input  wire d,
    output reg  q
);

    always @(posedge clk) begin
        if (rst)
            q <= 1'b0;      
        else if (en)
            q <= d;         
        else
            q <= q;        
    end

endmodule
